`timescale 1ns / 1ps
module name(clk,row,line);
    input clk;
    output [15:0] row;   //行输出
    output [3:0] line;   //列输出
    reg [3:0] count = 'd0; //控制哪一列被选中
    reg [9:0] num = 'd0;  //计数
    reg [2:0] S = 'd0;    //控制显示哪个汉字
    reg [3:0] line = 16'b1111111111111110; //列信号，在此初始化为选中第一列
    reg [15:0] row = 16'b0100000000001000; //行信号，在此初始化为第一个汉字在led上的第一列亮的那几个位置。

    always @(posedge clk) begin
        num = num + 1'b1;
        if (num > 10'd1023)
            num = 10'd00000000;
        else if (num == 10'd1023) begin //控制汉字的显示时间
            if (S == 4'd010) begin
                S = 3'b000;
            end else begin
                S = S + 1'b1;
            end
        end else begin
            S = S;
        end
    end

    always @(posedge clk) begin
        if (count < 4'd15) begin
            line = 3'b111; // 将所有列关闭，确保每次只有一列被选中。
            count = count + 1'd1;
        end else begin
            count = 4'd0;
        end
        // 由于line只有3位，我们不能直接使用line[count] = 1'b0的方式来选通某一列
        // 需要根据count的值来决定哪一位被置为0
        case (count[3:0])
            4'd0: line = 4'b0000;
            4'd1: line = 4'b0001;
            4'd2: line = 4'b0010;
            4'd3: line = 4'b0011;
            4'd4: line = 4'b0100;
            4'd5: line = 4'b0101;
            4'd6: line = 4'b0110;
            4'd7: line = 4'b0111;
            4'd8: line = 4'b1000;
            4'd9: line = 4'b1001;
            4'd10: line = 4'b1010;
            4'd11: line = 4'b1011;
            4'd12: line = 4'b1100;
            4'd13: line = 4'b1101;
            4'd14: line = 4'b1110;
            4'd15: line = 4'b1111;
            default: line = 4'b111; // 其他情况下关闭所有列
        endcase
    end

    always @(posedge clk) begin
        if (S == 4'b000) begin //王  左边为第15位，右边为第0位，每一串数字为一竖行
            case (count)
                4'b0000: row = 16'b0000000000000000;
                4'b0001: row = 16'b0000000000000000;
                4'b0010: row = 16'b0111111111111100;
                4'b0011: row = 16'b0000000100000000;
                4'b0100: row = 16'b0000000100000000;
                4'b0101: row = 16'b0000000100000000;
                4'b0110: row = 16'b0000000100000000;
                4'b0111: row = 16'b0000000100000000;
                4'b1000: row = 16'b0011111111111000;
                4'b1001: row = 16'b0000000100000000;
                4'b1010: row = 16'b0000000100000000;
                4'b1011: row = 16'b0000000100000000;
                4'b1100: row = 16'b0000000100000000;
                4'b1101: row = 16'b0000000100000000;
                4'b1110: row = 16'b1111111111111111;
                4'b1111: row = 16'b0000000000000000;
                default: row = 16'b0;
            endcase
        end else if (S == 4'b001) begin //文
            case (count)
                4'b0000: row = 16'b0000001000000000;
                4'b0001: row = 16'b0000000100000000;
                4'b0010: row = 16'b0000000100000000;
                4'b0011: row = 16'b1111111111111110;
                4'b0100: row = 16'b0001000000010000;
                4'b0101: row = 16'b0001000000010000;
                4'b0110: row = 16'b0000100000100000;
                4'b0111: row = 16'b0000100000100000;
                4'b1000: row = 16'b0000010001000000;
                4'b1001: row = 16'b0000001010000000;
                4'b1010: row = 16'b0000000100000000;
                4'b1011: row = 16'b0000001010000000;
                4'b1100: row = 16'b0000010001000000;
                4'b1101: row = 16'b0000100000100000;
                4'b1110: row = 16'b0011000000011000;
                4'b1111: row = 16'b1100000000000110;
                default: row = 16'b0;
            endcase
        end else if (S == 4'b010) begin //海
            case (count)
                4'b0000: row = 16'b0000000100000000;
                4'b0001: row = 16'b0010000100000000;
                4'b0010: row = 16'b0001000111111100;
                4'b0011: row = 16'b0001001000000000;
                4'b0100: row = 16'b1000010111111000;
                4'b0101: row = 16'b0100000100001000;
                4'b0110: row = 16'b0100100101001000;
                4'b0111: row = 16'b0000100100101000;
                4'b1000: row = 16'b0001011111111110;
                4'b1001: row = 16'b0001000100001000;
                4'b1010: row = 16'b1110001001001000;
                4'b1011: row = 16'b0010001000101000;
                4'b1100: row = 16'b0010001111111100;
                4'b1101: row = 16'b0010000000001000;
                4'b1110: row = 16'b0010000001010000;
                4'b1111: row = 16'b0000000000100000;
                default: row = 16'b0;
            endcase
        end else begin //什么都不显示
            case (count)
                4'b0000: row = 16'b0;
                4'b0001: row = 16'b0;
                4'b0010: row = 16'b0;
                4'b0011: row = 16'b0;
                4'b0100: row = 16'b0;
                4'b0101: row = 16'b0;
                4'b0110: row = 16'b0;
                4'b0111: row = 16'b0;
                4'b1000: row = 16'b0;
                4'b1001: row = 16'b0;
                4'b1010: row = 16'b0;
                4'b1011: row = 16'b0;
                4'b1100: row = 16'b0;
                4'b1101: row = 16'b0;
                4'b1110: row = 16'b0;
                4'b1111: row = 16'b0;
                default: row = 16'b0;
            endcase
        end
    end
endmodule